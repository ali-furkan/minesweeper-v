module main

import gg

fn main() {
	mut app := new_app()

	app.gg.run()
}
