module main

fn main() {
	mut app := new_app()

	app.gg.run()
}
